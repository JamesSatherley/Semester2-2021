library IEEE;
use IEEE.std_logic_1164.all;

entity Seven_seg is
	port ( x : in unsigned( 3 downto 0);
		seg : out std_logic_vector( 6 downto 0) );
end entity Seven_seg;


architecture comb of First is

begin

end architecture comb;
